logic a;
logic b;
always @ (posedge clk ) begin
  a <= b;
  end
